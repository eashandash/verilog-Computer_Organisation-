module csa64(s,c0,a,b,c);
    output  [63:0]s,c0;
    wire [63:0]s,c0;
    input [63:0]a,b,c;
    assign s=a^b^c;
    assign c0[0]=0;
	assign c0[1]=(a[0]&b[0])|(b[0]&c[0])|(c[0]&a[0]);
	assign c0[2]=(a[1]&b[1])|(b[1]&c[1])|(c[1]&a[1]);
	assign c0[3]=(a[2]&b[2])|(b[2]&c[2])|(c[2]&a[2]);
	assign c0[4]=(a[3]&b[3])|(b[3]&c[3])|(c[3]&a[3]);
	assign c0[5]=(a[4]&b[4])|(b[4]&c[4])|(c[4]&a[4]);
	assign c0[6]=(a[5]&b[5])|(b[5]&c[5])|(c[5]&a[5]);
	assign c0[7]=(a[6]&b[6])|(b[6]&c[6])|(c[6]&a[6]);
	assign c0[8]=(a[7]&b[7])|(b[7]&c[7])|(c[7]&a[7]);
	assign c0[9]=(a[8]&b[8])|(b[8]&c[8])|(c[8]&a[8]);
	assign c0[10]=(a[9]&b[9])|(b[9]&c[9])|(c[9]&a[9]);
	assign c0[11]=(a[10]&b[10])|(b[10]&c[10])|(c[10]&a[10]);
	assign c0[12]=(a[11]&b[11])|(b[11]&c[11])|(c[11]&a[11]);
	assign c0[13]=(a[12]&b[12])|(b[12]&c[12])|(c[12]&a[12]);
	assign c0[14]=(a[13]&b[13])|(b[13]&c[13])|(c[13]&a[13]);
	assign c0[15]=(a[14]&b[14])|(b[14]&c[14])|(c[14]&a[14]);
	assign c0[16]=(a[15]&b[15])|(b[15]&c[15])|(c[15]&a[15]);
	assign c0[17]=(a[16]&b[16])|(b[16]&c[16])|(c[16]&a[16]);
	assign c0[18]=(a[17]&b[17])|(b[17]&c[17])|(c[17]&a[17]);
	assign c0[19]=(a[18]&b[18])|(b[18]&c[18])|(c[18]&a[18]);
	assign c0[20]=(a[19]&b[19])|(b[19]&c[19])|(c[19]&a[19]);
	assign c0[21]=(a[20]&b[20])|(b[20]&c[20])|(c[20]&a[20]);
	assign c0[22]=(a[21]&b[21])|(b[21]&c[21])|(c[21]&a[21]);
	assign c0[23]=(a[22]&b[22])|(b[22]&c[22])|(c[22]&a[22]);
	assign c0[24]=(a[23]&b[23])|(b[23]&c[23])|(c[23]&a[23]);
	assign c0[25]=(a[24]&b[24])|(b[24]&c[24])|(c[24]&a[24]);
	assign c0[26]=(a[25]&b[25])|(b[25]&c[25])|(c[25]&a[25]);
	assign c0[27]=(a[26]&b[26])|(b[26]&c[26])|(c[26]&a[26]);
	assign c0[28]=(a[27]&b[27])|(b[27]&c[27])|(c[27]&a[27]);
	assign c0[29]=(a[28]&b[28])|(b[28]&c[28])|(c[28]&a[28]);
	assign c0[30]=(a[29]&b[29])|(b[29]&c[29])|(c[29]&a[29]);
	assign c0[31]=(a[30]&b[30])|(b[30]&c[30])|(c[30]&a[30]);
	assign c0[32]=(a[31]&b[31])|(b[31]&c[31])|(c[31]&a[31]);
	assign c0[33]=(a[32]&b[32])|(b[32]&c[32])|(c[32]&a[32]);
	assign c0[34]=(a[33]&b[33])|(b[33]&c[33])|(c[33]&a[33]);
	assign c0[35]=(a[34]&b[34])|(b[34]&c[34])|(c[34]&a[34]);
	assign c0[36]=(a[35]&b[35])|(b[35]&c[35])|(c[35]&a[35]);
	assign c0[37]=(a[36]&b[36])|(b[36]&c[36])|(c[36]&a[36]);
	assign c0[38]=(a[37]&b[37])|(b[37]&c[37])|(c[37]&a[37]);
	assign c0[39]=(a[38]&b[38])|(b[38]&c[38])|(c[38]&a[38]);
	assign c0[40]=(a[39]&b[39])|(b[39]&c[39])|(c[39]&a[39]);
	assign c0[41]=(a[40]&b[40])|(b[40]&c[40])|(c[40]&a[40]);
	assign c0[42]=(a[41]&b[41])|(b[41]&c[41])|(c[41]&a[41]);
	assign c0[43]=(a[42]&b[42])|(b[42]&c[42])|(c[42]&a[42]);
	assign c0[44]=(a[43]&b[43])|(b[43]&c[43])|(c[43]&a[43]);
	assign c0[45]=(a[44]&b[44])|(b[44]&c[44])|(c[44]&a[44]);
	assign c0[46]=(a[45]&b[45])|(b[45]&c[45])|(c[45]&a[45]);
	assign c0[47]=(a[46]&b[46])|(b[46]&c[46])|(c[46]&a[46]);
	assign c0[48]=(a[47]&b[47])|(b[47]&c[47])|(c[47]&a[47]);
	assign c0[49]=(a[48]&b[48])|(b[48]&c[48])|(c[48]&a[48]);
	assign c0[50]=(a[49]&b[49])|(b[49]&c[49])|(c[49]&a[49]);
	assign c0[51]=(a[50]&b[50])|(b[50]&c[50])|(c[50]&a[50]);
	assign c0[52]=(a[51]&b[51])|(b[51]&c[51])|(c[51]&a[51]);
	assign c0[53]=(a[52]&b[52])|(b[52]&c[52])|(c[52]&a[52]);
	assign c0[54]=(a[53]&b[53])|(b[53]&c[53])|(c[53]&a[53]);
	assign c0[55]=(a[54]&b[54])|(b[54]&c[54])|(c[54]&a[54]);
	assign c0[56]=(a[55]&b[55])|(b[55]&c[55])|(c[55]&a[55]);
	assign c0[57]=(a[56]&b[56])|(b[56]&c[56])|(c[56]&a[56]);
	assign c0[58]=(a[57]&b[57])|(b[57]&c[57])|(c[57]&a[57]);
	assign c0[59]=(a[58]&b[58])|(b[58]&c[58])|(c[58]&a[58]);
	assign c0[60]=(a[59]&b[59])|(b[59]&c[59])|(c[59]&a[59]);
	assign c0[61]=(a[60]&b[60])|(b[60]&c[60])|(c[60]&a[60]);
	assign c0[62]=(a[61]&b[61])|(b[61]&c[61])|(c[61]&a[61]);
	assign c0[63]=(a[62]&b[62])|(b[62]&c[62])|(c[62]&a[62]);




endmodule
