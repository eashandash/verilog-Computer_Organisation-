module ALU_tb();

reg [31:0]a2,a3,a4,a5,a6;
reg [31:0]b2,b3,b4,b5,b6,out1,out2;
wire [63:0]out3,out4,out5,out6;
//reg [4:0]opcode;
wire [63:0]OUT,L11,L12,L13,L21;


//exp^3
//taylor series till first 6 terms\

//term 2,3,4,5,6
//ALU t1(a2,b2,0111,out2);
ALU t2(a3,b3,0111,out3);
ALU t3(a4,b4,0111,out4);
ALU t4(a5,b5,0111,out5);
ALU t5(a6,b6,0111,out6);

//level 1
ALU l11(out1,out2,0101,L11);
ALU l12(out3[31:0],out4[31:0],0101,L12);
ALU l13(out5[31:0],out6[31:0],0101,L13);

//level 2
ALU l21(L11[31:0],L12[31:0],0101,L21);

//level 3
ALU l31(L13[31:0],L21[31:0],0101,OUT);

initial
begin
	out1=32'b00111111100000000000000000000000; 		//1
	out2=32'b01000000010000000000000000000000;		//3

	a3=32'b01000001000100000000000000000000;		//9
	b3=32'b00111111000000000000000000000000;		//0.5

	a4=32'b01000001110110000000000000000000;		//27
	b4=32'b00111110001010101010101010101011;       // 1/3!

	a5=32'b01000010101000100000000000000000;		//81
	b5=32'b00111101001010101010101010101011;	   // 1/4!

	a6=32'b01000011011100110000000000000000;		//243
	b6=32'b00111100000010001000100010001001;	   // 1/5!
end	

initial	
begin
$monitor("exp(3)=%b\n",OUT[31:0]);
end 	

endmodule // ALU_tb

