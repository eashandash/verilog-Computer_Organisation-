module imemory(addr, d_in, rd, wr, d_out);

   input [4:0]addr;
   input [31:0]d_in;
   input rd, wr;
   output [31:0]d_out;
   reg [31:0]d_out;

   reg [16:0]mem[16:0];
   



   initial
     begin
   	mem[0]=32'b0000_0000_0001_0010 ;
	mem[1]=32'b0010_0010_0011_0010 ;
	mem[2]=32'b0100_0010_0101_0010 ;
	mem[3]=32'b0110_0110_0111_0010 ;
	mem[4]=32'b1000_1000_1001_0010 ;
	mem[5]=32'b1010_1010_1011_0010 ;
	mem[6]=32'b1100_1100_1101_0010 ;
	mem[7]=32'b1110_1110_1111_0010 ;
	mem[8]=32'b0000_0000_0010_0010 ;	
	mem[9]=32'b0100_0100_0110_0010 ;	
	mem[10]=32'b1000_1000_1010_0010 ;	
	mem[11]=32'b1100_1100_1110_0010 ;	
	mem[12]=32'b0000_0000_0100_0010 ;
	mem[13]=32'b1000_1000_1100_0010 ;
	mem[14]=32'b0000_0000_1000_0010 ;

    end   
   










   always @ (*)
     begin

	if(rd == 1'b1)
	  begin
	     d_out <= mem[addr];
	  end
	

	else if(wr == 1'b1)
	  begin
	     mem[addr] <= d_in;
	  end
     end   
   
endmodule







module dmemory(addr, d_in, rd, wr, d_out);
   input[4:0] addr;
   input [31:0] d_in;
   input rd, wr;
   output [31:0] d_out;
   reg [31:0] d_out;
   reg [16:0]mem[31:0];
 
   

   initial
     begin
	mem[0]=32'b00111111100000000000000000000000;
	mem[1]=32'b01000001000100000000000000000000;
	mem[2]=32'b01000010001000100000000000000000;
	mem[3]=32'b01000010111100110000000000000000;
	mem[4]=32'b01000011100010001011000000000000;
	mem[5]=32'b01000011111101100000100110011010;
	mem[6]=32'b01000100001110001000011100110011;
	mem[7]=32'b01000100011011010100000000011101;
	mem[8]=32'b01000100100001010111010000010000;	
	mem[9]=32'b01000100100001010111010000010000;	
	mem[10]=32'b01000100011100000011011101010001;
	mem[11]=32'b01000100010001001000101001011001;
	mem[12]=32'b01000100000100110110011111000011;
	mem[13]=32'b01000011110011000001100110000100;
	mem[14]=32'b01000011100000110011010011111010;
	mem[15]=32'b01000011000111010111001011000101;	
     end
        
   




   always @ (*)
     begin

	if(rd == 1'b1)
	  begin
	     d_out = mem[addr];
	  end

	if(wr == 1'b1)
	  begin
	     mem[addr] = d_in;
	  end
     end

endmodule

