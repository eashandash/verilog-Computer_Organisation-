module wtm32(a,b,p,clk);
input [31:0]a,b;
input clk;
output [63:0]p;
wire [63:0]w1,w2,w3,w4,w5,w6,w7,w8,w9,w10,w11,w12,w13,w14,w15,w16,w17,w18,w19,w20,w21,w22,w23,w24,w25,w26,w27,w28,w29,w30,w31,w32;
wire  [63:0]wx1,wx2,wx3,wx4,wx5,wx6,wx7,wx8,wx9,wx10,wx11,wx12,wx13,wx14,wx15,wx16,wx17,wx18,wx19,wx20,wx21,wx22,wx23,wx24,wx25,wx26,wx27,wx28,wx29,wx30,wx31,wx32;
wire [63:0]s1,s2,s3,s4,s5,s6,s7,s8,s9,s10,s11,s12,s13,s14,s15,s16,s17,s18,s19,s20;
wire [63:0]k1,k2,k3,k4,k5,k6,k7,k8,k9,k10,k11,k12,k13,k14;
wire [63:0]l1,l2,l3,l4,l5,l6,l7,l8,l9,l10;
wire [63:0]m1,m2,m3,m4,m5,m6,qx1,qx2,px1,qx3,qx4,qx5,qx6,qx7,qx8,qx9,qx10,px2,px3,px4,px5;
wire [63:0]n1,n2,n3,n4;
wire q5,q4,q3,q6,q7,q8,q9;
wire [63:0]p1,p2,o1,o2,q1,q2,op1,op2,op3,op4,op5,op6,op7,op8;
//pp1
assign w1[0]= (a[0] & b[0]);
assign w1[1]= (a[0] & b[1]);
assign w1[2]= (a[0] & b[2]);
assign w1[3]= (a[0] & b[3]);
assign w1[4]= (a[0] & b[4]);
assign w1[5]= (a[0] & b[5]);
assign w1[6]= (a[0] & b[6]);
assign w1[7]= (a[0] & b[7]);
assign w1[8]= (a[0] & b[8]);
assign w1[9]= (a[0] & b[9]);
assign w1[10]= (a[0] & b[10]);
assign w1[11]= (a[0] & b[11]);
assign w1[12]= (a[0] & b[12]);
assign w1[13]= (a[0] & b[13]);
assign w1[14]= (a[0] & b[14]);
assign w1[15]= (a[0] & b[15]);
assign w1[16]= (a[0] & b[16]);
assign w1[17]= (a[0] & b[17]);
assign w1[18]= (a[0] & b[18]);
assign w1[19]= (a[0] & b[19]);
assign w1[20]= (a[0] & b[20]);
assign w1[21]= (a[0] & b[21]);
assign w1[22]= (a[0] & b[22]);
assign w1[23]= (a[0] & b[23]);
assign w1[24]= (a[0] & b[24]);
assign w1[25]= (a[0] & b[25]);
assign w1[26]= (a[0] & b[26]);
assign w1[27]= (a[0] & b[27]);
assign w1[28]= (a[0] & b[28]);
assign w1[29]= (a[0] & b[29]);
assign w1[30]= (a[0] & b[30]);
assign w1[31]= (a[0] & b[31]);
assign w1[63:32]= 0;
//pp2
assign w2[0]= 0 ;
assign w2[1]= (a[1] & b[0]);
assign w2[2]= (a[1] & b[1]);
assign w2[3]= (a[1] & b[2]);
assign w2[4]= (a[1] & b[3]);
assign w2[5]= (a[1] & b[4]);
assign w2[6]= (a[1] & b[5]);
assign w2[7]= (a[1] & b[6]);
assign w2[8]= (a[1] & b[7]);
assign w2[9]= (a[1] & b[8]);
assign w2[10]= (a[1] & b[9]);
assign w2[11]= (a[1] & b[10]);
assign w2[12]= (a[1] & b[11]);
assign w2[13]= (a[1] & b[12]);
assign w2[14]= (a[1] & b[13]);
assign w2[15]= (a[1] & b[14]);
assign w2[16]= (a[1] & b[15]);
assign w2[17]= (a[1] & b[16]);
assign w2[18]= (a[1] & b[17]);
assign w2[19]= (a[1] & b[18]);
assign w2[20]= (a[1] & b[19]);
assign w2[21]= (a[1] & b[20]);
assign w2[22]= (a[1] & b[21]);
assign w2[23]= (a[1] & b[22]);
assign w2[24]= (a[1] & b[23]);
assign w2[25]= (a[1] & b[24]);
assign w2[26]= (a[1] & b[25]);
assign w2[27]= (a[1] & b[26]);
assign w2[28]= (a[1] & b[27]);
assign w2[29]= (a[1] & b[28]);
assign w2[30]= (a[1] & b[29]);
assign w2[31]= (a[1] & b[30]);
assign w2[32]= (a[1] & b[31]);
assign w2[63:33]= 0 ;
//pp3
assign w3[0]= 0 ;
assign w3[1]= 0 ;
assign w3[2]= (a[2] & b[0]);
assign w3[3]= (a[2] & b[1]);
assign w3[4]= (a[2] & b[2]);
assign w3[5]= (a[2] & b[3]);
assign w3[6]= (a[2] & b[4]);
assign w3[7]= (a[2] & b[5]);
assign w3[8]= (a[2] & b[6]);
assign w3[9]= (a[2] & b[7]);
assign w3[10]= (a[2] & b[8]);
assign w3[11]= (a[2] & b[9]);
assign w3[12]= (a[2] & b[10]);
assign w3[13]= (a[2] & b[11]);
assign w3[14]= (a[2] & b[12]);
assign w3[15]= (a[2] & b[13]);
assign w3[16]= (a[2] & b[14]);
assign w3[17]= (a[2] & b[15]);
assign w3[18]= (a[2] & b[16]);
assign w3[19]= (a[2] & b[17]);
assign w3[20]= (a[2] & b[18]);
assign w3[21]= (a[2] & b[19]);
assign w3[22]= (a[2] & b[20]);
assign w3[23]= (a[2] & b[21]);
assign w3[24]= (a[2] & b[22]);
assign w3[25]= (a[2] & b[23]);
assign w3[26]= (a[2] & b[24]);
assign w3[27]= (a[2] & b[25]);
assign w3[28]= (a[2] & b[26]);
assign w3[29]= (a[2] & b[27]);
assign w3[30]= (a[2] & b[28]);
assign w3[31]= (a[2] & b[29]);
assign w3[32]= (a[2] & b[30]);
assign w3[33]= (a[2] & b[31]);
assign w3[63:34]= 0 ;
//pp4
assign w4[0]= 0 ;
assign w4[1]= 0 ;
assign w4[2]= 0 ;
assign w4[3]= (a[3] & b[0]);
assign w4[4]= (a[3] & b[1]);
assign w4[5]= (a[3] & b[2]);
assign w4[6]= (a[3] & b[3]);
assign w4[7]= (a[3] & b[4]);
assign w4[8]= (a[3] & b[5]);
assign w4[9]= (a[3] & b[6]);
assign w4[10]= (a[3] & b[7]);
assign w4[11]= (a[3] & b[8]);
assign w4[12]= (a[3] & b[9]);
assign w4[13]= (a[3] & b[10]);
assign w4[14]= (a[3] & b[11]);
assign w4[15]= (a[3] & b[12]);
assign w4[16]= (a[3] & b[13]);
assign w4[17]= (a[3] & b[14]);
assign w4[18]= (a[3] & b[15]);
assign w4[19]= (a[3] & b[16]);
assign w4[20]= (a[3] & b[17]);
assign w4[21]= (a[3] & b[18]);
assign w4[22]= (a[3] & b[19]);
assign w4[23]= (a[3] & b[20]);
assign w4[24]= (a[3] & b[21]);
assign w4[25]= (a[3] & b[22]);
assign w4[26]= (a[3] & b[23]);
assign w4[27]= (a[3] & b[24]);
assign w4[28]= (a[3] & b[25]);
assign w4[29]= (a[3] & b[26]);
assign w4[30]= (a[3] & b[27]);
assign w4[31]= (a[3] & b[28]);
assign w4[32]= (a[3] & b[29]);
assign w4[33]= (a[3] & b[30]);
assign w4[34]= (a[3] & b[31]);
assign w4[63:35]= 0 ;
//pp5
assign w5[3:0]= 0 ;
assign w5[4]= (a[4] & b[0]);
assign w5[5]= (a[4] & b[1]);
assign w5[6]= (a[4] & b[2]);
assign w5[7]= (a[4] & b[3]);
assign w5[8]= (a[4] & b[4]);
assign w5[9]= (a[4] & b[5]);
assign w5[10]= (a[4] & b[6]);
assign w5[11]= (a[4] & b[7]);
assign w5[12]= (a[4] & b[8]);
assign w5[13]= (a[4] & b[9]);
assign w5[14]= (a[4] & b[10]);
assign w5[15]= (a[4] & b[11]);
assign w5[16]= (a[4] & b[12]);
assign w5[17]= (a[4] & b[13]);
assign w5[18]= (a[4] & b[14]);
assign w5[19]= (a[4] & b[15]);
assign w5[20]= (a[4] & b[16]);
assign w5[21]= (a[4] & b[17]);
assign w5[22]= (a[4] & b[18]);
assign w5[23]= (a[4] & b[19]);
assign w5[24]= (a[4] & b[20]);
assign w5[25]= (a[4] & b[21]);
assign w5[26]= (a[4] & b[22]);
assign w5[27]= (a[4] & b[23]);
assign w5[28]= (a[4] & b[24]);
assign w5[29]= (a[4] & b[25]);
assign w5[30]= (a[4] & b[26]);
assign w5[31]= (a[4] & b[27]);
assign w5[32]= (a[4] & b[28]);
assign w5[33]= (a[4] & b[29]);
assign w5[34]= (a[4] & b[30]);
assign w5[35]= (a[4] & b[31]);
assign w5[63:36]= 0 ;
//pp6
assign w6[4:0]= 0 ;
assign w6[5]= (a[5] & b[0]);
assign w6[6]= (a[5] & b[1]);
assign w6[7]= (a[5] & b[2]);
assign w6[8]= (a[5] & b[3]);
assign w6[9]= (a[5] & b[4]);
assign w6[10]= (a[5] & b[5]);
assign w6[11]= (a[5] & b[6]);
assign w6[12]= (a[5] & b[7]);
assign w6[13]= (a[5] & b[8]);
assign w6[14]= (a[5] & b[9]);
assign w6[15]= (a[5] & b[10]);
assign w6[16]= (a[5] & b[11]);
assign w6[17]= (a[5] & b[12]);
assign w6[18]= (a[5] & b[13]);
assign w6[19]= (a[5] & b[14]);
assign w6[20]= (a[5] & b[15]);
assign w6[21]= (a[5] & b[16]);
assign w6[22]= (a[5] & b[17]);
assign w6[23]= (a[5] & b[18]);
assign w6[24]= (a[5] & b[19]);
assign w6[25]= (a[5] & b[20]);
assign w6[26]= (a[5] & b[21]);
assign w6[27]= (a[5] & b[22]);
assign w6[28]= (a[5] & b[23]);
assign w6[29]= (a[5] & b[24]);
assign w6[30]= (a[5] & b[25]);
assign w6[31]= (a[5] & b[26]);
assign w6[32]= (a[5] & b[27]);
assign w6[33]= (a[5] & b[28]);
assign w6[34]= (a[5] & b[29]);
assign w6[35]= (a[5] & b[30]);
assign w6[36]= (a[5] & b[31]);
assign w6[63:37]= 0 ;
//pp7
assign w7[5:0]= 0 ;
assign w7[6]= (a[6] & b[0]);
assign w7[7]= (a[6] & b[1]);
assign w7[8]= (a[6] & b[2]);
assign w7[9]= (a[6] & b[3]);
assign w7[10]= (a[6] & b[4]);
assign w7[11]= (a[6] & b[5]);
assign w7[12]= (a[6] & b[6]);
assign w7[13]= (a[6] & b[7]);
assign w7[14]= (a[6] & b[8]);
assign w7[15]= (a[6] & b[9]);
assign w7[16]= (a[6] & b[10]);
assign w7[17]= (a[6] & b[11]);
assign w7[18]= (a[6] & b[12]);
assign w7[19]= (a[6] & b[13]);
assign w7[20]= (a[6] & b[14]);
assign w7[21]= (a[6] & b[15]);
assign w7[22]= (a[6] & b[16]);
assign w7[23]= (a[6] & b[17]);
assign w7[24]= (a[6] & b[18]);
assign w7[25]= (a[6] & b[19]);
assign w7[26]= (a[6] & b[20]);
assign w7[27]= (a[6] & b[21]);
assign w7[28]= (a[6] & b[22]);
assign w7[29]= (a[6] & b[23]);
assign w7[30]= (a[6] & b[24]);
assign w7[31]= (a[6] & b[25]);
assign w7[32]= (a[6] & b[26]);
assign w7[33]= (a[6] & b[27]);
assign w7[34]= (a[6] & b[28]);
assign w7[35]= (a[6] & b[29]);
assign w7[36]= (a[6] & b[30]);
assign w7[37]= (a[6] & b[31]);
assign w7[63:38]= 0 ;
//pp8
assign w8[6:0]= 0 ;
assign w8[7]= (a[7] & b[0]);
assign w8[8]= (a[7] & b[1]);
assign w8[9]= (a[7] & b[2]);
assign w8[10]= (a[7] & b[3]);
assign w8[11]= (a[7] & b[4]);
assign w8[12]= (a[7] & b[5]);
assign w8[13]= (a[7] & b[6]);
assign w8[14]= (a[7] & b[7]);
assign w8[15]= (a[7] & b[8]);
assign w8[16]= (a[7] & b[9]);
assign w8[17]= (a[7] & b[10]);
assign w8[18]= (a[7] & b[11]);
assign w8[19]= (a[7] & b[12]);
assign w8[20]= (a[7] & b[13]);
assign w8[21]= (a[7] & b[14]);
assign w8[22]= (a[7] & b[15]);
assign w8[23]= (a[7] & b[16]);
assign w8[24]= (a[7] & b[17]);
assign w8[25]= (a[7] & b[18]);
assign w8[26]= (a[7] & b[19]);
assign w8[27]= (a[7] & b[20]);
assign w8[28]= (a[7] & b[21]);
assign w8[29]= (a[7] & b[22]);
assign w8[30]= (a[7] & b[23]);
assign w8[31]= (a[7] & b[24]);
assign w8[32]= (a[7] & b[25]);
assign w8[33]= (a[7] & b[26]);
assign w8[34]= (a[7] & b[27]);
assign w8[35]= (a[7] & b[28]);
assign w8[36]= (a[7] & b[29]);
assign w8[37]= (a[7] & b[30]);
assign w8[38]= (a[7] & b[31]);
assign w8[63:39]= 0 ;
//pp9
assign w9[7:0]= 0 ;
assign w9[8]= (a[8] & b[0]);
assign w9[9]= (a[8] & b[1]);
assign w9[10]= (a[8] & b[2]);
assign w9[11]= (a[8] & b[3]);
assign w9[12]= (a[8] & b[4]);
assign w9[13]= (a[8] & b[5]);
assign w9[14]= (a[8] & b[6]);
assign w9[15]= (a[8] & b[7]);
assign w9[16]= (a[8] & b[8]);
assign w9[17]= (a[8] & b[9]);
assign w9[18]= (a[8] & b[10]);
assign w9[19]= (a[8] & b[11]);
assign w9[20]= (a[8] & b[12]);
assign w9[21]= (a[8] & b[13]);
assign w9[22]= (a[8] & b[14]);
assign w9[23]= (a[8] & b[15]);
assign w9[24]= (a[8] & b[16]);
assign w9[25]= (a[8] & b[17]);
assign w9[26]= (a[8] & b[18]);
assign w9[27]= (a[8] & b[19]);
assign w9[28]= (a[8] & b[20]);
assign w9[29]= (a[8] & b[21]);
assign w9[30]= (a[8] & b[22]);
assign w9[31]= (a[8] & b[23]);
assign w9[32]= (a[8] & b[24]);
assign w9[33]= (a[8] & b[25]);
assign w9[34]= (a[8] & b[26]);
assign w9[35]= (a[8] & b[27]);
assign w9[36]= (a[8] & b[28]);
assign w9[37]= (a[8] & b[29]);
assign w9[38]= (a[8] & b[30]);
assign w9[39]= (a[8] & b[31]);
assign w9[63:40]= 0 ;
//pp10
assign w10[8:0]= 0 ;
assign w10[9]= (a[9] & b[0]);
assign w10[10]= (a[9] & b[1]);
assign w10[11]= (a[9] & b[2]);
assign w10[12]= (a[9] & b[3]);
assign w10[13]= (a[9] & b[4]);
assign w10[14]= (a[9] & b[5]);
assign w10[15]= (a[9] & b[6]);
assign w10[16]= (a[9] & b[7]);
assign w10[17]= (a[9] & b[8]);
assign w10[18]= (a[9] & b[9]);
assign w10[19]= (a[9] & b[10]);
assign w10[20]= (a[9] & b[11]);
assign w10[21]= (a[9] & b[12]);
assign w10[22]= (a[9] & b[13]);
assign w10[23]= (a[9] & b[14]);
assign w10[24]= (a[9] & b[15]);
assign w10[25]= (a[9] & b[16]);
assign w10[26]= (a[9] & b[17]);
assign w10[27]= (a[9] & b[18]);
assign w10[28]= (a[9] & b[19]);
assign w10[29]= (a[9] & b[20]);
assign w10[30]= (a[9] & b[21]);
assign w10[31]= (a[9] & b[22]);
assign w10[32]= (a[9] & b[23]);
assign w10[33]= (a[9] & b[24]);
assign w10[34]= (a[9] & b[25]);
assign w10[35]= (a[9] & b[26]);
assign w10[36]= (a[9] & b[27]);
assign w10[37]= (a[9] & b[28]);
assign w10[38]= (a[9] & b[29]);
assign w10[39]= (a[9] & b[30]);
assign w10[40]= (a[9] & b[31]);
assign w10[63:41]= 0 ;
//pp11
assign w11[9:0]= 0 ;
assign w11[10]= (a[10] & b[0]);
assign w11[11]= (a[10] & b[1]);
assign w11[12]= (a[10] & b[2]);
assign w11[13]= (a[10] & b[3]);
assign w11[14]= (a[10] & b[4]);
assign w11[15]= (a[10] & b[5]);
assign w11[16]= (a[10] & b[6]);
assign w11[17]= (a[10] & b[7]);
assign w11[18]= (a[10] & b[8]);
assign w11[19]= (a[10] & b[9]);
assign w11[20]= (a[10] & b[10]);
assign w11[21]= (a[10] & b[11]);
assign w11[22]= (a[10] & b[12]);
assign w11[23]= (a[10] & b[13]);
assign w11[24]= (a[10] & b[14]);
assign w11[25]= (a[10] & b[15]);
assign w11[26]= (a[10] & b[16]);
assign w11[27]= (a[10] & b[17]);
assign w11[28]= (a[10] & b[18]);
assign w11[29]= (a[10] & b[19]);
assign w11[30]= (a[10] & b[20]);
assign w11[31]= (a[10] & b[21]);
assign w11[32]= (a[10] & b[22]);
assign w11[33]= (a[10] & b[23]);
assign w11[34]= (a[10] & b[24]);
assign w11[35]= (a[10] & b[25]);
assign w11[36]= (a[10] & b[26]);
assign w11[37]= (a[10] & b[27]);
assign w11[38]= (a[10] & b[28]);
assign w11[39]= (a[10] & b[29]);
assign w11[40]= (a[10] & b[30]);
assign w11[41]= (a[10] & b[31]);
assign w11[63:42]= 0 ;
//pp12
assign w12[10:0]= 0 ;
assign w12[11]= (a[11] & b[0]);
assign w12[12]= (a[11] & b[1]);
assign w12[13]= (a[11] & b[2]);
assign w12[14]= (a[11] & b[3]);
assign w12[15]= (a[11] & b[4]);
assign w12[16]= (a[11] & b[5]);
assign w12[17]= (a[11] & b[6]);
assign w12[18]= (a[11] & b[7]);
assign w12[19]= (a[11] & b[8]);
assign w12[20]= (a[11] & b[9]);
assign w12[21]= (a[11] & b[10]);
assign w12[22]= (a[11] & b[11]);
assign w12[23]= (a[11] & b[12]);
assign w12[24]= (a[11] & b[13]);
assign w12[25]= (a[11] & b[14]);
assign w12[26]= (a[11] & b[15]);
assign w12[27]= (a[11] & b[16]);
assign w12[28]= (a[11] & b[17]);
assign w12[29]= (a[11] & b[18]);
assign w12[30]= (a[11] & b[19]);
assign w12[31]= (a[11] & b[20]);
assign w12[32]= (a[11] & b[21]);
assign w12[33]= (a[11] & b[22]);
assign w12[34]= (a[11] & b[23]);
assign w12[35]= (a[11] & b[24]);
assign w12[36]= (a[11] & b[25]);
assign w12[37]= (a[11] & b[26]);
assign w12[38]= (a[11] & b[27]);
assign w12[39]= (a[11] & b[28]);
assign w12[40]= (a[11] & b[29]);
assign w12[41]= (a[11] & b[30]);
assign w12[42]= (a[11] & b[31]);
assign w12[63:43]= 0 ;
//pp13
assign w13[11:0]= 0 ;
assign w13[12]= (a[12] & b[0]);
assign w13[13]= (a[12] & b[1]);
assign w13[14]= (a[12] & b[2]);
assign w13[15]= (a[12] & b[3]);
assign w13[16]= (a[12] & b[4]);
assign w13[17]= (a[12] & b[5]);
assign w13[18]= (a[12] & b[6]);
assign w13[19]= (a[12] & b[7]);
assign w13[20]= (a[12] & b[8]);
assign w13[21]= (a[12] & b[9]);
assign w13[22]= (a[12] & b[10]);
assign w13[23]= (a[12] & b[11]);
assign w13[24]= (a[12] & b[12]);
assign w13[25]= (a[12] & b[13]);
assign w13[26]= (a[12] & b[14]);
assign w13[27]= (a[12] & b[15]);
assign w13[28]= (a[12] & b[16]);
assign w13[29]= (a[12] & b[17]);
assign w13[30]= (a[12] & b[18]);
assign w13[31]= (a[12] & b[19]);
assign w13[32]= (a[12] & b[20]);
assign w13[33]= (a[12] & b[21]);
assign w13[34]= (a[12] & b[22]);
assign w13[35]= (a[12] & b[23]);
assign w13[36]= (a[12] & b[24]);
assign w13[37]= (a[12] & b[25]);
assign w13[38]= (a[12] & b[26]);
assign w13[39]= (a[12] & b[27]);
assign w13[40]= (a[12] & b[28]);
assign w13[41]= (a[12] & b[29]);
assign w13[42]= (a[12] & b[30]);
assign w13[43]= (a[12] & b[31]);
assign w13[63:44]= 0 ;
//pp14
assign w14[12:0]= 0 ;
assign w14[13]= (a[13] & b[0]);
assign w14[14]= (a[13] & b[1]);
assign w14[15]= (a[13] & b[2]);
assign w14[16]= (a[13] & b[3]);
assign w14[17]= (a[13] & b[4]);
assign w14[18]= (a[13] & b[5]);
assign w14[19]= (a[13] & b[6]);
assign w14[20]= (a[13] & b[7]);
assign w14[21]= (a[13] & b[8]);
assign w14[22]= (a[13] & b[9]);
assign w14[23]= (a[13] & b[10]);
assign w14[24]= (a[13] & b[11]);
assign w14[25]= (a[13] & b[12]);
assign w14[26]= (a[13] & b[13]);
assign w14[27]= (a[13] & b[14]);
assign w14[28]= (a[13] & b[15]);
assign w14[29]= (a[13] & b[16]);
assign w14[30]= (a[13] & b[17]);
assign w14[31]= (a[13] & b[18]);
assign w14[32]= (a[13] & b[19]);
assign w14[33]= (a[13] & b[20]);
assign w14[34]= (a[13] & b[21]);
assign w14[35]= (a[13] & b[22]);
assign w14[36]= (a[13] & b[23]);
assign w14[37]= (a[13] & b[24]);
assign w14[38]= (a[13] & b[25]);
assign w14[39]= (a[13] & b[26]);
assign w14[40]= (a[13] & b[27]);
assign w14[41]= (a[13] & b[28]);
assign w14[42]= (a[13] & b[29]);
assign w14[43]= (a[13] & b[30]);
assign w14[44]= (a[13] & b[31]);
assign w14[63:45]= 0 ;
//pp15
assign w15[13:0]= 0 ;
assign w15[14]= (a[14] & b[0]);
assign w15[15]= (a[14] & b[1]);
assign w15[16]= (a[14] & b[2]);
assign w15[17]= (a[14] & b[3]);
assign w15[18]= (a[14] & b[4]);
assign w15[19]= (a[14] & b[5]);
assign w15[20]= (a[14] & b[6]);
assign w15[21]= (a[14] & b[7]);
assign w15[22]= (a[14] & b[8]);
assign w15[23]= (a[14] & b[9]);
assign w15[24]= (a[14] & b[10]);
assign w15[25]= (a[14] & b[11]);
assign w15[26]= (a[14] & b[12]);
assign w15[27]= (a[14] & b[13]);
assign w15[28]= (a[14] & b[14]);
assign w15[29]= (a[14] & b[15]);
assign w15[30]= (a[14] & b[16]);
assign w15[31]= (a[14] & b[17]);
assign w15[32]= (a[14] & b[18]);
assign w15[33]= (a[14] & b[19]);
assign w15[34]= (a[14] & b[20]);
assign w15[35]= (a[14] & b[21]);
assign w15[36]= (a[14] & b[22]);
assign w15[37]= (a[14] & b[23]);
assign w15[38]= (a[14] & b[24]);
assign w15[39]= (a[14] & b[25]);
assign w15[40]= (a[14] & b[26]);
assign w15[41]= (a[14] & b[27]);
assign w15[42]= (a[14] & b[28]);
assign w15[43]= (a[14] & b[29]);
assign w15[44]= (a[14] & b[30]);
assign w15[45]= (a[14] & b[31]);
assign w15[63:46]= 0 ;
//pp16
assign w16[14:0]= 0 ;
assign w16[15]= (a[15] & b[0]);
assign w16[16]= (a[15] & b[1]);
assign w16[17]= (a[15] & b[2]);
assign w16[18]= (a[15] & b[3]);
assign w16[19]= (a[15] & b[4]);
assign w16[20]= (a[15] & b[5]);
assign w16[21]= (a[15] & b[6]);
assign w16[22]= (a[15] & b[7]);
assign w16[23]= (a[15] & b[8]);
assign w16[24]= (a[15] & b[9]);
assign w16[25]= (a[15] & b[10]);
assign w16[26]= (a[15] & b[11]);
assign w16[27]= (a[15] & b[12]);
assign w16[28]= (a[15] & b[13]);
assign w16[29]= (a[15] & b[14]);
assign w16[30]= (a[15] & b[15]);
assign w16[31]= (a[15] & b[16]);
assign w16[32]= (a[15] & b[17]);
assign w16[33]= (a[15] & b[18]);
assign w16[34]= (a[15] & b[19]);
assign w16[35]= (a[15] & b[20]);
assign w16[36]= (a[15] & b[21]);
assign w16[37]= (a[15] & b[22]);
assign w16[38]= (a[15] & b[23]);
assign w16[39]= (a[15] & b[24]);
assign w16[40]= (a[15] & b[25]);
assign w16[41]= (a[15] & b[26]);
assign w16[42]= (a[15] & b[27]);
assign w16[43]= (a[15] & b[28]);
assign w16[44]= (a[15] & b[29]);
assign w16[45]= (a[15] & b[30]);
assign w16[46]= (a[15] & b[31]);
assign w16[63:47]= 0 ;
//pp17
assign w17[15:0]= 0 ;
assign w17[16]= (a[16] & b[0]);
assign w17[17]= (a[16] & b[1]);
assign w17[18]= (a[16] & b[2]);
assign w17[19]= (a[16] & b[3]);
assign w17[20]= (a[16] & b[4]);
assign w17[21]= (a[16] & b[5]);
assign w17[22]= (a[16] & b[6]);
assign w17[23]= (a[16] & b[7]);
assign w17[24]= (a[16] & b[8]);
assign w17[25]= (a[16] & b[9]);
assign w17[26]= (a[16] & b[10]);
assign w17[27]= (a[16] & b[11]);
assign w17[28]= (a[16] & b[12]);
assign w17[29]= (a[16] & b[13]);
assign w17[30]= (a[16] & b[14]);
assign w17[31]= (a[16] & b[15]);
assign w17[32]= (a[16] & b[16]);
assign w17[33]= (a[16] & b[17]);
assign w17[34]= (a[16] & b[18]);
assign w17[35]= (a[16] & b[19]);
assign w17[36]= (a[16] & b[20]);
assign w17[37]= (a[16] & b[21]);
assign w17[38]= (a[16] & b[22]);
assign w17[39]= (a[16] & b[23]);
assign w17[40]= (a[16] & b[24]);
assign w17[41]= (a[16] & b[25]);
assign w17[42]= (a[16] & b[26]);
assign w17[43]= (a[16] & b[27]);
assign w17[44]= (a[16] & b[28]);
assign w17[45]= (a[16] & b[29]);
assign w17[46]= (a[16] & b[30]);
assign w17[47]= (a[16] & b[31]);
assign w17[63:48]= 0 ;
//pp18
assign w18[16:0]= 0 ;
assign w18[17]= (a[17] & b[0]);
assign w18[18]= (a[17] & b[1]);
assign w18[19]= (a[17] & b[2]);
assign w18[20]= (a[17] & b[3]);
assign w18[21]= (a[17] & b[4]);
assign w18[22]= (a[17] & b[5]);
assign w18[23]= (a[17] & b[6]);
assign w18[24]= (a[17] & b[7]);
assign w18[25]= (a[17] & b[8]);
assign w18[26]= (a[17] & b[9]);
assign w18[27]= (a[17] & b[10]);
assign w18[28]= (a[17] & b[11]);
assign w18[29]= (a[17] & b[12]);
assign w18[30]= (a[17] & b[13]);
assign w18[31]= (a[17] & b[14]);
assign w18[32]= (a[17] & b[15]);
assign w18[33]= (a[17] & b[16]);
assign w18[34]= (a[17] & b[17]);
assign w18[35]= (a[17] & b[18]);
assign w18[36]= (a[17] & b[19]);
assign w18[37]= (a[17] & b[20]);
assign w18[38]= (a[17] & b[21]);
assign w18[39]= (a[17] & b[22]);
assign w18[40]= (a[17] & b[23]);
assign w18[41]= (a[17] & b[24]);
assign w18[42]= (a[17] & b[25]);
assign w18[43]= (a[17] & b[26]);
assign w18[44]= (a[17] & b[27]);
assign w18[45]= (a[17] & b[28]);
assign w18[46]= (a[17] & b[29]);
assign w18[47]= (a[17] & b[30]);
assign w18[48]= (a[17] & b[31]);
assign w18[63:49]= 0 ;
//pp19
assign w19[17:0]= 0 ;
assign w19[18]= (a[18] & b[0]);
assign w19[19]= (a[18] & b[1]);
assign w19[20]= (a[18] & b[2]);
assign w19[21]= (a[18] & b[3]);
assign w19[22]= (a[18] & b[4]);
assign w19[23]= (a[18] & b[5]);
assign w19[24]= (a[18] & b[6]);
assign w19[25]= (a[18] & b[7]);
assign w19[26]= (a[18] & b[8]);
assign w19[27]= (a[18] & b[9]);
assign w19[28]= (a[18] & b[10]);
assign w19[29]= (a[18] & b[11]);
assign w19[30]= (a[18] & b[12]);
assign w19[31]= (a[18] & b[13]);
assign w19[32]= (a[18] & b[14]);
assign w19[33]= (a[18] & b[15]);
assign w19[34]= (a[18] & b[16]);
assign w19[35]= (a[18] & b[17]);
assign w19[36]= (a[18] & b[18]);
assign w19[37]= (a[18] & b[19]);
assign w19[38]= (a[18] & b[20]);
assign w19[39]= (a[18] & b[21]);
assign w19[40]= (a[18] & b[22]);
assign w19[41]= (a[18] & b[23]);
assign w19[42]= (a[18] & b[24]);
assign w19[43]= (a[18] & b[25]);
assign w19[44]= (a[18] & b[26]);
assign w19[45]= (a[18] & b[27]);
assign w19[46]= (a[18] & b[28]);
assign w19[47]= (a[18] & b[29]);
assign w19[48]= (a[18] & b[30]);
assign w19[49]= (a[18] & b[31]);
assign w19[63:50]= 0 ;
//pp20
assign w20[18:0]= 0 ;
assign w20[19]= (a[19] & b[0]);
assign w20[20]= (a[19] & b[1]);
assign w20[21]= (a[19] & b[2]);
assign w20[22]= (a[19] & b[3]);
assign w20[23]= (a[19] & b[4]);
assign w20[24]= (a[19] & b[5]);
assign w20[25]= (a[19] & b[6]);
assign w20[26]= (a[19] & b[7]);
assign w20[27]= (a[19] & b[8]);
assign w20[28]= (a[19] & b[9]);
assign w20[29]= (a[19] & b[10]);
assign w20[30]= (a[19] & b[11]);
assign w20[31]= (a[19] & b[12]);
assign w20[32]= (a[19] & b[13]);
assign w20[33]= (a[19] & b[14]);
assign w20[34]= (a[19] & b[15]);
assign w20[35]= (a[19] & b[16]);
assign w20[36]= (a[19] & b[17]);
assign w20[37]= (a[19] & b[18]);
assign w20[38]= (a[19] & b[19]);
assign w20[39]= (a[19] & b[20]);
assign w20[40]= (a[19] & b[21]);
assign w20[41]= (a[19] & b[22]);
assign w20[42]= (a[19] & b[23]);
assign w20[43]= (a[19] & b[24]);
assign w20[44]= (a[19] & b[25]);
assign w20[45]= (a[19] & b[26]);
assign w20[46]= (a[19] & b[27]);
assign w20[47]= (a[19] & b[28]);
assign w20[48]= (a[19] & b[29]);
assign w20[49]= (a[19] & b[30]);
assign w20[50]= (a[19] & b[31]);
assign w20[63:51]= 0 ;
//pp21
assign w21[19:0]= 0 ;
assign w21[20]= (a[20] & b[0]);
assign w21[21]= (a[20] & b[1]);
assign w21[22]= (a[20] & b[2]);
assign w21[23]= (a[20] & b[3]);
assign w21[24]= (a[20] & b[4]);
assign w21[25]= (a[20] & b[5]);
assign w21[26]= (a[20] & b[6]);
assign w21[27]= (a[20] & b[7]);
assign w21[28]= (a[20] & b[8]);
assign w21[29]= (a[20] & b[9]);
assign w21[30]= (a[20] & b[10]);
assign w21[31]= (a[20] & b[11]);
assign w21[32]= (a[20] & b[12]);
assign w21[33]= (a[20] & b[13]);
assign w21[34]= (a[20] & b[14]);
assign w21[35]= (a[20] & b[15]);
assign w21[36]= (a[20] & b[16]);
assign w21[37]= (a[20] & b[17]);
assign w21[38]= (a[20] & b[18]);
assign w21[39]= (a[20] & b[19]);
assign w21[40]= (a[20] & b[20]);
assign w21[41]= (a[20] & b[21]);
assign w21[42]= (a[20] & b[22]);
assign w21[43]= (a[20] & b[23]);
assign w21[44]= (a[20] & b[24]);
assign w21[45]= (a[20] & b[25]);
assign w21[46]= (a[20] & b[26]);
assign w21[47]= (a[20] & b[27]);
assign w21[48]= (a[20] & b[28]);
assign w21[49]= (a[20] & b[29]);
assign w21[50]= (a[20] & b[30]);
assign w21[51]= (a[20] & b[31]);
assign w21[63:52]= 0 ;
//pp22
assign w22[20:0]= 0 ;
assign w22[21]= (a[21] & b[0]);
assign w22[22]= (a[21] & b[1]);
assign w22[23]= (a[21] & b[2]);
assign w22[24]= (a[21] & b[3]);
assign w22[25]= (a[21] & b[4]);
assign w22[26]= (a[21] & b[5]);
assign w22[27]= (a[21] & b[6]);
assign w22[28]= (a[21] & b[7]);
assign w22[29]= (a[21] & b[8]);
assign w22[30]= (a[21] & b[9]);
assign w22[31]= (a[21] & b[10]);
assign w22[32]= (a[21] & b[11]);
assign w22[33]= (a[21] & b[12]);
assign w22[34]= (a[21] & b[13]);
assign w22[35]= (a[21] & b[14]);
assign w22[36]= (a[21] & b[15]);
assign w22[37]= (a[21] & b[16]);
assign w22[38]= (a[21] & b[17]);
assign w22[39]= (a[21] & b[18]);
assign w22[40]= (a[21] & b[19]);
assign w22[41]= (a[21] & b[20]);
assign w22[42]= (a[21] & b[21]);
assign w22[43]= (a[21] & b[22]);
assign w22[44]= (a[21] & b[23]);
assign w22[45]= (a[21] & b[24]);
assign w22[46]= (a[21] & b[25]);
assign w22[47]= (a[21] & b[26]);
assign w22[48]= (a[21] & b[27]);
assign w22[49]= (a[21] & b[28]);
assign w22[50]= (a[21] & b[29]);
assign w22[51]= (a[21] & b[30]);
assign w22[52]= (a[21] & b[31]);
assign w22[63:53]= 0 ;
//pp23
assign w23[21:0]= 0 ;
assign w23[22]= (a[22] & b[0]);
assign w23[23]= (a[22] & b[1]);
assign w23[24]= (a[22] & b[2]);
assign w23[25]= (a[22] & b[3]);
assign w23[26]= (a[22] & b[4]);
assign w23[27]= (a[22] & b[5]);
assign w23[28]= (a[22] & b[6]);
assign w23[29]= (a[22] & b[7]);
assign w23[30]= (a[22] & b[8]);
assign w23[31]= (a[22] & b[9]);
assign w23[32]= (a[22] & b[10]);
assign w23[33]= (a[22] & b[11]);
assign w23[34]= (a[22] & b[12]);
assign w23[35]= (a[22] & b[13]);
assign w23[36]= (a[22] & b[14]);
assign w23[37]= (a[22] & b[15]);
assign w23[38]= (a[22] & b[16]);
assign w23[39]= (a[22] & b[17]);
assign w23[40]= (a[22] & b[18]);
assign w23[41]= (a[22] & b[19]);
assign w23[42]= (a[22] & b[20]);
assign w23[43]= (a[22] & b[21]);
assign w23[44]= (a[22] & b[22]);
assign w23[45]= (a[22] & b[23]);
assign w23[46]= (a[22] & b[24]);
assign w23[47]= (a[22] & b[25]);
assign w23[48]= (a[22] & b[26]);
assign w23[49]= (a[22] & b[27]);
assign w23[50]= (a[22] & b[28]);
assign w23[51]= (a[22] & b[29]);
assign w23[52]= (a[22] & b[30]);
assign w23[53]= (a[22] & b[31]);
assign w23[63:54]= 0 ;
//pp24
assign w24[22:0]= 0 ;
assign w24[23]= (a[23] & b[0]);
assign w24[24]= (a[23] & b[1]);
assign w24[25]= (a[23] & b[2]);
assign w24[26]= (a[23] & b[3]);
assign w24[27]= (a[23] & b[4]);
assign w24[28]= (a[23] & b[5]);
assign w24[29]= (a[23] & b[6]);
assign w24[30]= (a[23] & b[7]);
assign w24[31]= (a[23] & b[8]);
assign w24[32]= (a[23] & b[9]);
assign w24[33]= (a[23] & b[10]);
assign w24[34]= (a[23] & b[11]);
assign w24[35]= (a[23] & b[12]);
assign w24[36]= (a[23] & b[13]);
assign w24[37]= (a[23] & b[14]);
assign w24[38]= (a[23] & b[15]);
assign w24[39]= (a[23] & b[16]);
assign w24[40]= (a[23] & b[17]);
assign w24[41]= (a[23] & b[18]);
assign w24[42]= (a[23] & b[19]);
assign w24[43]= (a[23] & b[20]);
assign w24[44]= (a[23] & b[21]);
assign w24[45]= (a[23] & b[22]);
assign w24[46]= (a[23] & b[23]);
assign w24[47]= (a[23] & b[24]);
assign w24[48]= (a[23] & b[25]);
assign w24[49]= (a[23] & b[26]);
assign w24[50]= (a[23] & b[27]);
assign w24[51]= (a[23] & b[28]);
assign w24[52]= (a[23] & b[29]);
assign w24[53]= (a[23] & b[30]);
assign w24[54]= (a[23] & b[31]);
assign w24[63:55]= 0 ;
//pp25
assign w25[23:0]= 0 ;
assign w25[24]= (a[24] & b[0]);
assign w25[25]= (a[24] & b[1]);
assign w25[26]= (a[24] & b[2]);
assign w25[27]= (a[24] & b[3]);
assign w25[28]= (a[24] & b[4]);
assign w25[29]= (a[24] & b[5]);
assign w25[30]= (a[24] & b[6]);
assign w25[31]= (a[24] & b[7]);
assign w25[32]= (a[24] & b[8]);
assign w25[33]= (a[24] & b[9]);
assign w25[34]= (a[24] & b[10]);
assign w25[35]= (a[24] & b[11]);
assign w25[36]= (a[24] & b[12]);
assign w25[37]= (a[24] & b[13]);
assign w25[38]= (a[24] & b[14]);
assign w25[39]= (a[24] & b[15]);
assign w25[40]= (a[24] & b[16]);
assign w25[41]= (a[24] & b[17]);
assign w25[42]= (a[24] & b[18]);
assign w25[43]= (a[24] & b[19]);
assign w25[44]= (a[24] & b[20]);
assign w25[45]= (a[24] & b[21]);
assign w25[46]= (a[24] & b[22]);
assign w25[47]= (a[24] & b[23]);
assign w25[48]= (a[24] & b[24]);
assign w25[49]= (a[24] & b[25]);
assign w25[50]= (a[24] & b[26]);
assign w25[51]= (a[24] & b[27]);
assign w25[52]= (a[24] & b[28]);
assign w25[53]= (a[24] & b[29]);
assign w25[54]= (a[24] & b[30]);
assign w25[55]= (a[24] & b[31]);
assign w25[63:56]= 0 ;
//pp26
assign w26[24:0]= 0 ;
assign w26[25]= (a[25] & b[0]);
assign w26[26]= (a[25] & b[1]);
assign w26[27]= (a[25] & b[2]);
assign w26[28]= (a[25] & b[3]);
assign w26[29]= (a[25] & b[4]);
assign w26[30]= (a[25] & b[5]);
assign w26[31]= (a[25] & b[6]);
assign w26[32]= (a[25] & b[7]);
assign w26[33]= (a[25] & b[8]);
assign w26[34]= (a[25] & b[9]);
assign w26[35]= (a[25] & b[10]);
assign w26[36]= (a[25] & b[11]);
assign w26[37]= (a[25] & b[12]);
assign w26[38]= (a[25] & b[13]);
assign w26[39]= (a[25] & b[14]);
assign w26[40]= (a[25] & b[15]);
assign w26[41]= (a[25] & b[16]);
assign w26[42]= (a[25] & b[17]);
assign w26[43]= (a[25] & b[18]);
assign w26[44]= (a[25] & b[19]);
assign w26[45]= (a[25] & b[20]);
assign w26[46]= (a[25] & b[21]);
assign w26[47]= (a[25] & b[22]);
assign w26[48]= (a[25] & b[23]);
assign w26[49]= (a[25] & b[24]);
assign w26[50]= (a[25] & b[25]);
assign w26[51]= (a[25] & b[26]);
assign w26[52]= (a[25] & b[27]);
assign w26[53]= (a[25] & b[28]);
assign w26[54]= (a[25] & b[29]);
assign w26[55]= (a[25] & b[30]);
assign w26[56]= (a[25] & b[31]);
assign w26[63:57]= 0 ;
//pp27
assign w27[25:0]= 0 ;
assign w27[26]= (a[26] & b[0]);
assign w27[27]= (a[26] & b[1]);
assign w27[28]= (a[26] & b[2]);
assign w27[29]= (a[26] & b[3]);
assign w27[30]= (a[26] & b[4]);
assign w27[31]= (a[26] & b[5]);
assign w27[32]= (a[26] & b[6]);
assign w27[33]= (a[26] & b[7]);
assign w27[34]= (a[26] & b[8]);
assign w27[35]= (a[26] & b[9]);
assign w27[36]= (a[26] & b[10]);
assign w27[37]= (a[26] & b[11]);
assign w27[38]= (a[26] & b[12]);
assign w27[39]= (a[26] & b[13]);
assign w27[40]= (a[26] & b[14]);
assign w27[41]= (a[26] & b[15]);
assign w27[42]= (a[26] & b[16]);
assign w27[43]= (a[26] & b[17]);
assign w27[44]= (a[26] & b[18]);
assign w27[45]= (a[26] & b[19]);
assign w27[46]= (a[26] & b[20]);
assign w27[47]= (a[26] & b[21]);
assign w27[48]= (a[26] & b[22]);
assign w27[49]= (a[26] & b[23]);
assign w27[50]= (a[26] & b[24]);
assign w27[51]= (a[26] & b[25]);
assign w27[52]= (a[26] & b[26]);
assign w27[53]= (a[26] & b[27]);
assign w27[54]= (a[26] & b[28]);
assign w27[55]= (a[26] & b[29]);
assign w27[56]= (a[26] & b[30]);
assign w27[57]= (a[26] & b[31]);
assign w27[63:58]= 0 ;
//pp28
assign w28[26:0]= 0 ;
assign w28[27]= (a[27] & b[0]);
assign w28[28]= (a[27] & b[1]);
assign w28[29]= (a[27] & b[2]);
assign w28[30]= (a[27] & b[3]);
assign w28[31]= (a[27] & b[4]);
assign w28[32]= (a[27] & b[5]);
assign w28[33]= (a[27] & b[6]);
assign w28[34]= (a[27] & b[7]);
assign w28[35]= (a[27] & b[8]);
assign w28[36]= (a[27] & b[9]);
assign w28[37]= (a[27] & b[10]);
assign w28[38]= (a[27] & b[11]);
assign w28[39]= (a[27] & b[12]);
assign w28[40]= (a[27] & b[13]);
assign w28[41]= (a[27] & b[14]);
assign w28[42]= (a[27] & b[15]);
assign w28[43]= (a[27] & b[16]);
assign w28[44]= (a[27] & b[17]);
assign w28[45]= (a[27] & b[18]);
assign w28[46]= (a[27] & b[19]);
assign w28[47]= (a[27] & b[20]);
assign w28[48]= (a[27] & b[21]);
assign w28[49]= (a[27] & b[22]);
assign w28[50]= (a[27] & b[23]);
assign w28[51]= (a[27] & b[24]);
assign w28[52]= (a[27] & b[25]);
assign w28[53]= (a[27] & b[26]);
assign w28[54]= (a[27] & b[27]);
assign w28[55]= (a[27] & b[28]);
assign w28[56]= (a[27] & b[29]);
assign w28[57]= (a[27] & b[30]);
assign w28[58]= (a[27] & b[31]);
assign w28[63:59]= 0 ;
//pp29
assign w29[27:0]= 0 ;
assign w29[28]= (a[28] & b[0]);
assign w29[29]= (a[28] & b[1]);
assign w29[30]= (a[28] & b[2]);
assign w29[31]= (a[28] & b[3]);
assign w29[32]= (a[28] & b[4]);
assign w29[33]= (a[28] & b[5]);
assign w29[34]= (a[28] & b[6]);
assign w29[35]= (a[28] & b[7]);
assign w29[36]= (a[28] & b[8]);
assign w29[37]= (a[28] & b[9]);
assign w29[38]= (a[28] & b[10]);
assign w29[39]= (a[28] & b[11]);
assign w29[40]= (a[28] & b[12]);
assign w29[41]= (a[28] & b[13]);
assign w29[42]= (a[28] & b[14]);
assign w29[43]= (a[28] & b[15]);
assign w29[44]= (a[28] & b[16]);
assign w29[45]= (a[28] & b[17]);
assign w29[46]= (a[28] & b[18]);
assign w29[47]= (a[28] & b[19]);
assign w29[48]= (a[28] & b[20]);
assign w29[49]= (a[28] & b[21]);
assign w29[50]= (a[28] & b[22]);
assign w29[51]= (a[28] & b[23]);
assign w29[52]= (a[28] & b[24]);
assign w29[53]= (a[28] & b[25]);
assign w29[54]= (a[28] & b[26]);
assign w29[55]= (a[28] & b[27]);
assign w29[56]= (a[28] & b[28]);
assign w29[57]= (a[28] & b[29]);
assign w29[58]= (a[28] & b[30]);
assign w29[59]= (a[28] & b[31]);
assign w29[63:60]= 0 ;
//pp30
assign w30[28:0]= 0 ;
assign w30[29]= (a[29] & b[0]);
assign w30[30]= (a[29] & b[1]);
assign w30[31]= (a[29] & b[2]);
assign w30[32]= (a[29] & b[3]);
assign w30[33]= (a[29] & b[4]);
assign w30[34]= (a[29] & b[5]);
assign w30[35]= (a[29] & b[6]);
assign w30[36]= (a[29] & b[7]);
assign w30[37]= (a[29] & b[8]);
assign w30[38]= (a[29] & b[9]);
assign w30[39]= (a[29] & b[10]);
assign w30[40]= (a[29] & b[11]);
assign w30[41]= (a[29] & b[12]);
assign w30[42]= (a[29] & b[13]);
assign w30[43]= (a[29] & b[14]);
assign w30[44]= (a[29] & b[15]);
assign w30[45]= (a[29] & b[16]);
assign w30[46]= (a[29] & b[17]);
assign w30[47]= (a[29] & b[18]);
assign w30[48]= (a[29] & b[19]);
assign w30[49]= (a[29] & b[20]);
assign w30[50]= (a[29] & b[21]);
assign w30[51]= (a[29] & b[22]);
assign w30[52]= (a[29] & b[23]);
assign w30[53]= (a[29] & b[24]);
assign w30[54]= (a[29] & b[25]);
assign w30[55]= (a[29] & b[26]);
assign w30[56]= (a[29] & b[27]);
assign w30[57]= (a[29] & b[28]);
assign w30[58]= (a[29] & b[29]);
assign w30[59]= (a[29] & b[30]);
assign w30[60]= (a[29] & b[31]);
assign w30[63:61]= 0 ;
//pp31
assign w31[29:0]= 0 ;
assign w31[30]= (a[30] & b[0]);
assign w31[31]= (a[30] & b[1]);
assign w31[32]= (a[30] & b[2]);
assign w31[33]= (a[30] & b[3]);
assign w31[34]= (a[30] & b[4]);
assign w31[35]= (a[30] & b[5]);
assign w31[36]= (a[30] & b[6]);
assign w31[37]= (a[30] & b[7]);
assign w31[38]= (a[30] & b[8]);
assign w31[39]= (a[30] & b[9]);
assign w31[40]= (a[30] & b[10]);
assign w31[41]= (a[30] & b[11]);
assign w31[42]= (a[30] & b[12]);
assign w31[43]= (a[30] & b[13]);
assign w31[44]= (a[30] & b[14]);
assign w31[45]= (a[30] & b[15]);
assign w31[46]= (a[30] & b[16]);
assign w31[47]= (a[30] & b[17]);
assign w31[48]= (a[30] & b[18]);
assign w31[49]= (a[30] & b[19]);
assign w31[50]= (a[30] & b[20]);
assign w31[51]= (a[30] & b[21]);
assign w31[52]= (a[30] & b[22]);
assign w31[53]= (a[30] & b[23]);
assign w31[54]= (a[30] & b[24]);
assign w31[55]= (a[30] & b[25]);
assign w31[56]= (a[30] & b[26]);
assign w31[57]= (a[30] & b[27]);
assign w31[58]= (a[30] & b[28]);
assign w31[59]= (a[30] & b[29]);
assign w31[60]= (a[30] & b[30]);
assign w31[61]= (a[30] & b[31]);
assign w31[63:62]= 0 ;
//pp32
assign w32[30:0]= 0 ;
assign w32[31]= (a[31] & b[0]);
assign w32[32]= (a[31] & b[1]);
assign w32[33]= (a[31] & b[2]);
assign w32[34]= (a[31] & b[3]);
assign w32[35]= (a[31] & b[4]);
assign w32[36]= (a[31] & b[5]);
assign w32[37]= (a[31] & b[6]);
assign w32[38]= (a[31] & b[7]);
assign w32[39]= (a[31] & b[8]);
assign w32[40]= (a[31] & b[9]);
assign w32[41]= (a[31] & b[10]);
assign w32[42]= (a[31] & b[11]);
assign w32[43]= (a[31] & b[12]);
assign w32[44]= (a[31] & b[13]);
assign w32[45]= (a[31] & b[14]);
assign w32[46]= (a[31] & b[15]);
assign w32[47]= (a[31] & b[16]);
assign w32[48]= (a[31] & b[17]);
assign w32[49]= (a[31] & b[18]);
assign w32[50]= (a[31] & b[19]);
assign w32[51]= (a[31] & b[20]);
assign w32[52]= (a[31] & b[21]);
assign w32[53]= (a[31] & b[22]);
assign w32[54]= (a[31] & b[23]);
assign w32[55]= (a[31] & b[24]);
assign w32[56]= (a[31] & b[25]);
assign w32[57]= (a[31] & b[26]);
assign w32[58]= (a[31] & b[27]);
assign w32[59]= (a[31] & b[28]);
assign w32[60]= (a[31] & b[29]);
assign w32[61]= (a[31] & b[30]);
assign w32[62]= (a[31] & b[31]);
assign w32[63]= 0 ;
//passing pp to dff_64
dff_64 ff1(wx1,w1,clk);
dff_64 ff2(wx2,w2,clk);
dff_64 ff3(wx3,w3,clk);
dff_64 ff4(wx4,w4,clk);
dff_64 ff5(wx5,w5,clk);
dff_64 ff6(wx6,w6,clk);
dff_64 ff7(wx7,w7,clk);
dff_64 ff8(wx8,w8,clk);
dff_64 ff9(wx9,w9,clk);
dff_64 ff10(wx10,w10,clk);
dff_64 ff11(wx11,w11,clk);
dff_64 ff12(wx12,w12,clk);
dff_64 ff13(wx13,w13,clk);
dff_64 ff14(wx14,w14,clk);
dff_64 ff15(wx15,w15,clk);
dff_64 ff16(wx16,w16,clk);
dff_64 ff17(wx17,w17,clk);
dff_64 ff18(wx18,w18,clk);
dff_64 ff19(wx19,w19,clk);
dff_64 ff20(wx20,w20,clk);
dff_64 ff21(wx21,w21,clk);
dff_64 ff22(wx22,w22,clk);
dff_64 ff23(wx23,w23,clk);
dff_64 ff24(wx24,w24,clk);
dff_64 ff25(wx25,w25,clk);
dff_64 ff26(wx26,w26,clk);
dff_64 ff27(wx27,w27,clk);
dff_64 ff28(wx28,w28,clk);
dff_64 ff29(wx29,w29,clk);
dff_64 ff30(wx30,w30,clk);
dff_64 ff31(wx31,w31,clk);
dff_64 ff32(wx32,w32,clk);

//assign p=wx3;
//level 1 csa
csa a1(wx1,wx2,wx3,s1,s2,clk);
csa a2(wx4,wx5,wx6,s3,s4,clk);
csa a3(wx7,wx8,wx9,s5,s6,clk);
csa a4(wx10,wx11,wx12,s7,s8,clk);
csa a5(wx13,wx14,wx15,s9,s10,clk);
csa a6(wx16,wx17,wx18,s11,s12,clk);
csa a7(wx19,wx20,wx21,s13,s14,clk);
csa a8(wx22,wx23,wx24,s15,s16,clk);
csa a9(wx25,wx26,wx27,s17,s18,clk);
csa a10(wx28,wx29,wx30,s19,s20,clk);
dff_64 ff33(op1,wx31,clk);
dff_64 ff34(op2,wx32,clk);
//level 2 csa
csa b1(s1,s2,s3,k1,k2,clk);
csa b2(s4,s5,s6,k3,k4,clk);
csa b3(s7,s8,s9,k5,k6,clk);
csa b4(s10,s11,s12,k7,k8,clk);
csa b5(s13,s14,s15,k9,k10,clk);
csa b6(s16,s17,s18,k11,k12,clk);
csa b7(s19,s20,op1,k13,k14,clk);
dff_64 ff35(op3,op2,clk);
//level 3 csa
csa c1(k1,k2,k3,l1,l2,clk);
csa c2(k4,k5,k6,l3,l4,clk);
csa c3(k7,k8,k9,l5,l6,clk);
csa c4(k10,k11,k12,l7,l8,clk);
csa c5(k13,k14,op3,l9,l10,clk);
//level 4 csa
csa d1(l1,l2,l3,m1,m2,clk);
csa d2(l4,l5,l6,m3,m4,clk);
csa d3(l7,l8,l9,m5,m6,clk);
dff_64 ff36(op4,l10,clk);
//level 5 csa
csa e1(m1,m2,m3,n1,n2,clk);
csa e2(m4,m5,m6,n3,n4,clk);
dff_64 ff37(op5,op4,clk);
//level 6 csa
csa f1(n1,n2,n3,p1,p2,clk);
dff_64 ff38(op6,op5,clk);
dff_64 ff39(op7,n4,clk);
//level 7 csa
csa g1(p1,p2,op7,o1,o2,clk);
dff_64 ff40(op8,op6,clk);
//level 8
csa g2(o1,o2,op8,q1,q2,clk);
//assign p=q2;
pre32p y1(px1[31:0],q4,q1[31:0],q2[31:0],0,clk);
dff_32 ff43(qx1[63:32],q1[63:32],clk);
dff_32 ff44(qx2[63:32],q2[63:32],clk);
dff_32 ff47(qx3[63:32],qx1[63:32],clk);
dff_32 ff48(qx4[63:32],qx2[63:32],clk);


dff_32 ff51(qx5[63:32],qx3[63:32],clk);
dff_32 ff52(qx6[63:32],qx4[63:32],clk);

dff_32 ff55(qx7[63:32],qx5[63:32],clk);
dff_32 ff56(qx8[63:32],qx6[63:32],clk);

dff_32 ff59(qx9[63:32],qx7[63:32],clk);
dff_32 ff60(qx10[63:32],qx8[63:32],clk);

pre32p y2(p[63:32],q3,qx9[63:32],qx10[63:32],q4,clk);

dff_32 ff42(px2[31:0],px1[31:0],clk);
dff_32 ff46(px3[31:0],px2[31:0],clk);
dff_32 ff50(px4[31:0],px3[31:0],clk);
dff_32 ff54(px5[31:0],px4[31:0],clk);
dff_32 ff58(p[31:0],px5[31:0],clk);

endmodule


